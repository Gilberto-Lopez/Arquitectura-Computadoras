`timescale 1ns / 1ps
//Test Sumador de 32 bits con signo
module TestSumador;

	//Inputs
	reg [31:0] a;
	reg [31:0] b;
	//Outputs
	wire [31:0] Z;
	wire ovf;

	//Unit under test
	Sumador uut(
		.a(a),
		.b(b),
		.Z(Z),
		.ovf(ovf)
	);
	
	initial begin
		a = 32'b0;
		b = 32'b0;

		#100;

		a = 32'h0; b = 32'h0; //0+0
		#50;
		$display("Z = %b %b.%b, ovf = %b", Z[31], Z[30:10], Z[9:0], ovf);
		a = 32'h0; b = 32'h80000000; //0+(-0)
		#50;
		$display("Z = %b %b.%b, ovf = %b", Z[31], Z[30:10], Z[9:0], ovf);
		a = 32'h80000000; b = 32'h0; //-0+0
		#50;
		$display("Z = %b %b.%b, ovf = %b", Z[31], Z[30:10], Z[9:0], ovf);
		a = 32'h200; b = 32'h400; //.1 + 1
		#50;
		$display("Z = %b %b.%b, ovf = %b", Z[31], Z[30:10], Z[9:0], ovf);
		a = 32'h508; b = 32'h989680; //1.0100001 + 10011000100101.101
		#50;
		$display("Z = %b %b.%b, ovf = %b", Z[31], Z[30:10], Z[9:0], ovf);
		a = 32'hA8D99763; b = 32'hDE6D23E4; //-10100011011001100101.1101100011 + -101111001101101001000.11111001
		#50;
		$display("Z = %b %b.%b, ovf = %b", Z[31], Z[30:10], Z[9:0], ovf);
		a = 32'h28D99763; b = 32'h5E6D23E4; //10100011011001100101.1101100011 + 101111001101101001000.11111001
		#50;
		$display("Z = %b %b.%b, ovf = %b", Z[31], Z[30:10], Z[9:0], ovf);
		a = 32'hB2EF5901; b = 32'h35905D0E; //-11001011101111010110.0100000001 + 11010110010000010111.010000111
		#50;
		$display("Z = %b %b.%b, ovf = %b", Z[31], Z[30:10], Z[9:0], ovf);
		a = 32'h14C7DBC7; b = 32'h8DFAE342; //1010011000111110110.1111000111 + -110111111010111000.110100001
		#50;
		$display("Z = %b %b.%b, ovf = %b", Z[31], Z[30:10], Z[9:0], ovf);
		a = 32'h94C7DBC7; b = 32'hDFAE342; //-1010011000111110110.1111000111 + 110111111010111000.110100001
		#50;
		$display("Z = %b %b.%b, ovf = %b", Z[31], Z[30:10], Z[9:0], ovf);
	end

endmodule
